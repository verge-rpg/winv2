#define OBJECTS 30

#define NOTHING         1
#define VANISHING       2
#define HURTPLAYER      4
#define HURTENEMIES     8
#define OBSTRUCTABLE    16
#define EXPLOSIVE       32

#define DIR_UP          0
#define DIR_LEFT        270
#define DIR_DOWN        180
#define DIR_RIGHT       90
